-- Copyright (C) 2016  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 16.1.0 Build 196 10/24/2016 SJ Lite Edition
-- Created on Sat Oct 17 15:57:06 2020

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY HW6P2 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        A : IN STD_LOGIC := '0';
        B : IN STD_LOGIC := '0';
        C : IN STD_LOGIC := '0';
        D : IN STD_LOGIC := '0';
        PBGNT : IN STD_LOGIC := '0';
        MACK : IN STD_LOGIC := '0';
        CON : IN STD_LOGIC := '0';
        PBREQ : OUT STD_LOGIC;
        CMREQ : OUT STD_LOGIC;
        CE : OUT STD_LOGIC;
        CNTLD : OUT STD_LOGIC;
        CLD : OUT STD_LOGIC
    );
END HW6P2;

ARCHITECTURE BEHAVIOR OF HW6P2 IS
    TYPE type_fstate IS (state0,state4,state5,state1,state2,state3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,A,B,C,D,PBGNT,MACK,CON)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state0;
            PBREQ <= '0';
            CMREQ <= '0';
            CE <= '0';
            CNTLD <= '0';
            CLD <= '0';
        ELSE
            PBREQ <= '0';
            CMREQ <= '0';
            CE <= '0';
            CNTLD <= '0';
            CLD <= '0';
            CASE fstate IS
                WHEN state0 =>
                    IF (((((A = '1') AND (B = '1')) AND (C = '1')) AND (D = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF (((((A = '0') AND (B = '0')) AND (C = '0')) AND (D = '0'))) THEN
                        reg_fstate <= state0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state0;
                    END IF;
                WHEN state4 =>
                    IF ((CON = '1')) THEN
                        reg_fstate <= state5;
                    ELSIF ((CON = '0')) THEN
                        reg_fstate <= state0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    CLD <= '1';
                WHEN state5 =>
                    IF ((MACK = '1')) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    CMREQ <= '1';
                WHEN state1 =>
                    IF ((PBGNT = '1')) THEN
                        reg_fstate <= state2;
                    ELSIF ((PBGNT = '0')) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    PBREQ <= '1';
                WHEN state2 =>
                    IF ((MACK = '1')) THEN
                        reg_fstate <= state3;
                    ELSIF ((MACK = '0')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    CNTLD <= '1';

                    CMREQ <= '1';
                WHEN state3 =>
                    IF ((MACK = '1')) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    CE <= '1';
                WHEN OTHERS => 
                    PBREQ <= 'X';
                    CMREQ <= 'X';
                    CE <= 'X';
                    CNTLD <= 'X';
                    CLD <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
