LIBRARY altera_mf;USE
        altera_mf.altera_mf_components.all;
		  