// Copyright (C) 2016  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus Prime Version 16.1.0 Build 196 10/24/2016 SJ Lite Edition
// Created on Sat Oct 17 16:01:06 2020

// synthesis message_off 10175

`timescale 1ns/1ns

module HW6P2 (
    reset,clock,A,B,C,D,PBGNT,MACK,CON,
    PBREQ,CMREQ,CE,CNTLD,CLD);

    input reset;
    input clock;
    input A;
    input B;
    input C;
    input D;
    input PBGNT;
    input MACK;
    input CON;
    tri0 reset;
    tri0 A;
    tri0 B;
    tri0 C;
    tri0 D;
    tri0 PBGNT;
    tri0 MACK;
    tri0 CON;
    output PBREQ;
    output CMREQ;
    output CE;
    output CNTLD;
    output CLD;
    reg PBREQ;
    reg CMREQ;
    reg CE;
    reg CNTLD;
    reg CLD;
    reg [5:0] fstate;
    reg [5:0] reg_fstate;
    parameter state0=0,state4=1,state5=2,state1=3,state2=4,state3=5;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or A or B or C or D or PBGNT or MACK or CON)
    begin
        if (reset) begin
            reg_fstate <= state0;
            PBREQ <= 1'b0;
            CMREQ <= 1'b0;
            CE <= 1'b0;
            CNTLD <= 1'b0;
            CLD <= 1'b0;
        end
        else begin
            PBREQ <= 1'b0;
            CMREQ <= 1'b0;
            CE <= 1'b0;
            CNTLD <= 1'b0;
            CLD <= 1'b0;
            case (fstate)
                state0: begin
                    if (((((A == 1'b1) & (B == 1'b1)) & (C == 1'b1)) & (D == 1'b1)))
                        reg_fstate <= state1;
                    else if (((((A == 1'b0) & (B == 1'b0)) & (C == 1'b0)) & (D == 1'b0)))
                        reg_fstate <= state0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state0;
                end
                state4: begin
                    if ((CON == 1'b1))
                        reg_fstate <= state5;
                    else if ((CON == 1'b0))
                        reg_fstate <= state0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    CLD <= 1'b1;
                end
                state5: begin
                    if ((MACK == 1'b1))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    CMREQ <= 1'b1;
                end
                state1: begin
                    if ((PBGNT == 1'b1))
                        reg_fstate <= state2;
                    else if ((PBGNT == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    PBREQ <= 1'b1;
                end
                state2: begin
                    if ((MACK == 1'b1))
                        reg_fstate <= state3;
                    else if ((MACK == 1'b0))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    CNTLD <= 1'b1;

                    CMREQ <= 1'b1;
                end
                state3: begin
                    if ((MACK == 1'b1))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    CE <= 1'b1;
                end
                default: begin
                    PBREQ <= 1'bx;
                    CMREQ <= 1'bx;
                    CE <= 1'bx;
                    CNTLD <= 1'bx;
                    CLD <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // HW6P2
